CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 330 421 0 1 3
0 10
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89883e-315 0
0
6 74LS48
188 983 655 0 14 29
0 13 15 2 11 17 18 9 8 7
6 5 4 3 19
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 665 427 0 3 22
0 16 15 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3536 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 475 418 0 3 22
0 11 2 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4597 0 0
2
5.89883e-315 0
0
6 74112~
219 851 482 0 7 32
0 10 14 12 14 10 20 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
3835 0 0
2
5.89883e-315 0
0
6 74112~
219 591 608 0 7 32
0 10 16 12 16 10 21 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6A
-25 -64 -4 -56
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
3670 0 0
2
5.89883e-315 0
0
6 74112~
219 447 605 0 7 32
0 10 11 12 11 10 2 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 4 0
1 U
5616 0 0
2
5.89883e-315 0
0
6 74112~
219 330 628 0 7 32
0 10 22 12 23 10 24 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
9323 0 0
2
5.89883e-315 0
0
7 Pulser~
4 250 601 0 10 12
0 25 26 27 12 0 0 5 2 4
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
317 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 1116 456 0 18 19
10 3 4 5 6 7 8 9 28 29
1 1 1 1 0 0 1 2 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3108 0 0
2
5.89883e-315 5.26354e-315
0
36
6 0 2 0 0 8192 0 7 0 0 30 4
477 587
475 587
475 617
486 617
13 1 3 0 0 8320 0 2 10 0 0 3
1015 673
1095 673
1095 492
12 2 4 0 0 8320 0 2 10 0 0 3
1015 664
1101 664
1101 492
11 3 5 0 0 8320 0 2 10 0 0 3
1015 655
1107 655
1107 492
10 4 6 0 0 8320 0 2 10 0 0 3
1015 646
1113 646
1113 492
9 5 7 0 0 8320 0 2 10 0 0 3
1015 637
1119 637
1119 492
8 6 8 0 0 8320 0 2 10 0 0 3
1015 628
1125 628
1125 492
7 7 9 0 0 8320 0 2 10 0 0 3
1015 619
1131 619
1131 492
0 0 10 0 0 4096 0 0 0 21 14 2
376 504
376 707
0 0 10 0 0 0 0 0 0 21 13 2
511 504
511 707
0 0 10 0 0 0 0 0 0 21 12 2
667 504
667 706
0 5 10 0 0 8192 0 0 5 13 0 4
584 707
584 706
851 706
851 494
0 5 10 0 0 0 0 0 6 14 0 3
446 707
591 707
591 620
5 5 10 0 0 0 0 8 7 0 0 4
330 640
330 707
447 707
447 617
0 1 11 0 0 8192 0 0 4 16 0 4
401 617
389 617
389 409
451 409
4 2 11 0 0 0 0 7 7 0 0 6
423 587
401 587
401 617
395 617
395 569
423 569
3 3 12 0 0 12416 0 7 6 0 0 6
417 578
412 578
412 668
532 668
532 581
561 581
1 0 10 0 0 0 0 1 0 0 21 2
330 430
330 504
1 0 10 0 0 0 0 6 0 0 21 2
591 545
591 504
1 0 10 0 0 0 0 7 0 0 21 2
447 542
447 504
1 1 10 0 0 8320 0 5 8 0 0 4
851 419
851 504
330 504
330 565
7 1 13 0 0 12416 0 5 2 0 0 4
875 446
776 446
776 619
951 619
2 3 14 0 0 8320 0 5 3 0 0 3
827 446
827 427
686 427
2 4 14 0 0 4224 0 5 5 0 0 4
827 446
684 446
684 464
827 464
7 2 15 0 0 12416 0 6 2 0 0 4
615 572
658 572
658 628
951 628
7 2 15 0 0 0 0 6 3 0 0 4
615 572
618 572
618 436
641 436
4 2 16 0 0 8192 0 6 6 0 0 4
567 590
555 590
555 572
567 572
2 3 16 0 0 8320 0 6 4 0 0 4
567 572
555 572
555 418
496 418
7 4 11 0 0 12416 0 8 2 0 0 4
354 592
383 592
383 646
951 646
7 3 2 0 0 12416 0 7 2 0 0 4
471 569
486 569
486 637
951 637
7 2 2 0 0 0 0 7 4 0 0 4
471 569
441 569
441 427
451 427
7 2 11 0 0 0 0 8 7 0 0 4
354 592
416 592
416 569
423 569
3 4 12 0 0 128 0 8 9 0 0 2
300 601
280 601
3 3 12 0 0 16512 0 6 5 0 0 6
561 581
550 581
550 668
676 668
676 455
821 455
3 3 12 0 0 0 0 8 7 0 0 6
300 601
294 601
294 668
406 668
406 578
417 578
3 1 16 0 0 16 0 4 3 0 0 2
496 418
641 418
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
